
`ifndef CAPTURE_SV
`define CAPTURE_SV

`endif
